`ifndef BLOCK_0_VH
`define BLOCK_0_VH
`define BLOCK_0_REGISTER_0_BIT_FIELD_0_BIT_WIDTH 4
`define BLOCK_0_REGISTER_0_BIT_FIELD_0_BIT_MASK 4'hf
`define BLOCK_0_REGISTER_0_BIT_FIELD_0_BIT_OFFSET 0
`define BLOCK_0_REGISTER_0_BIT_FIELD_1_BIT_WIDTH 4
`define BLOCK_0_REGISTER_0_BIT_FIELD_1_BIT_MASK 4'hf
`define BLOCK_0_REGISTER_0_BIT_FIELD_1_BIT_OFFSET 4
`define BLOCK_0_REGISTER_0_BIT_FIELD_2_BIT_WIDTH 1
`define BLOCK_0_REGISTER_0_BIT_FIELD_2_BIT_MASK 1'h1
`define BLOCK_0_REGISTER_0_BIT_FIELD_2_BIT_OFFSET 8
`define BLOCK_0_REGISTER_0_BIT_FIELD_3_BIT_WIDTH 2
`define BLOCK_0_REGISTER_0_BIT_FIELD_3_BIT_MASK 2'h3
`define BLOCK_0_REGISTER_0_BIT_FIELD_3_BIT_OFFSET 9
`define BLOCK_0_REGISTER_0_BIT_FIELD_4_BIT_WIDTH 2
`define BLOCK_0_REGISTER_0_BIT_FIELD_4_BIT_MASK 2'h3
`define BLOCK_0_REGISTER_0_BIT_FIELD_4_BIT_OFFSET 11
`define BLOCK_0_REGISTER_0_BIT_FIELD_5_BIT_WIDTH 2
`define BLOCK_0_REGISTER_0_BIT_FIELD_5_BIT_MASK 2'h3
`define BLOCK_0_REGISTER_0_BIT_FIELD_5_BIT_OFFSET 13
`define BLOCK_0_REGISTER_0_BIT_FIELD_6_BIT_WIDTH 2
`define BLOCK_0_REGISTER_0_BIT_FIELD_6_BIT_MASK 2'h3
`define BLOCK_0_REGISTER_0_BIT_FIELD_6_BIT_OFFSET 15
`define BLOCK_0_REGISTER_0_BYTE_WIDTH 4
`define BLOCK_0_REGISTER_0_BYTE_SIZE 4
`define BLOCK_0_REGISTER_0_BYTE_OFFSET 8'h00
`define BLOCK_0_REGISTER_1_BIT_WIDTH 1
`define BLOCK_0_REGISTER_1_BIT_MASK 1'h1
`define BLOCK_0_REGISTER_1_BIT_OFFSET 0
`define BLOCK_0_REGISTER_1_FOO 1'h0
`define BLOCK_0_REGISTER_1_BAR 1'h1
`define BLOCK_0_REGISTER_1_BYTE_WIDTH 4
`define BLOCK_0_REGISTER_1_BYTE_SIZE 4
`define BLOCK_0_REGISTER_1_BYTE_OFFSET 8'h04
`define BLOCK_0_REGISTER_2_BIT_FIELD_0_BIT_WIDTH 4
`define BLOCK_0_REGISTER_2_BIT_FIELD_0_BIT_MASK 4'hf
`define BLOCK_0_REGISTER_2_BIT_FIELD_0_BIT_OFFSET 0
`define BLOCK_0_REGISTER_2_BIT_FIELD_1_BIT_WIDTH 8
`define BLOCK_0_REGISTER_2_BIT_FIELD_1_BIT_MASK 8'hff
`define BLOCK_0_REGISTER_2_BIT_FIELD_1_BIT_OFFSET 8
`define BLOCK_0_REGISTER_2_BIT_FIELD_2_BIT_WIDTH 4
`define BLOCK_0_REGISTER_2_BIT_FIELD_2_BIT_MASK 4'hf
`define BLOCK_0_REGISTER_2_BIT_FIELD_2_BIT_OFFSET 16
`define BLOCK_0_REGISTER_2_BIT_FIELD_3_BIT_WIDTH 4
`define BLOCK_0_REGISTER_2_BIT_FIELD_3_BIT_MASK 4'hf
`define BLOCK_0_REGISTER_2_BIT_FIELD_3_BIT_OFFSET 20
`define BLOCK_0_REGISTER_2_BYTE_WIDTH 4
`define BLOCK_0_REGISTER_2_BYTE_SIZE 4
`define BLOCK_0_REGISTER_2_BYTE_OFFSET 8'h08
`define BLOCK_0_REGISTER_3_BIT_FIELD_0_BIT_WIDTH 4
`define BLOCK_0_REGISTER_3_BIT_FIELD_0_BIT_MASK 4'hf
`define BLOCK_0_REGISTER_3_BIT_FIELD_0_BIT_OFFSET 0
`define BLOCK_0_REGISTER_3_BIT_FIELD_1_BIT_WIDTH 4
`define BLOCK_0_REGISTER_3_BIT_FIELD_1_BIT_MASK 4'hf
`define BLOCK_0_REGISTER_3_BIT_FIELD_1_BIT_OFFSET 4
`define BLOCK_0_REGISTER_3_BIT_FIELD_2_BIT_WIDTH 4
`define BLOCK_0_REGISTER_3_BIT_FIELD_2_BIT_MASK 4'hf
`define BLOCK_0_REGISTER_3_BIT_FIELD_2_BIT_OFFSET 8
`define BLOCK_0_REGISTER_3_BIT_FIELD_3_BIT_WIDTH 4
`define BLOCK_0_REGISTER_3_BIT_FIELD_3_BIT_MASK 4'hf
`define BLOCK_0_REGISTER_3_BIT_FIELD_3_BIT_OFFSET 16
`define BLOCK_0_REGISTER_3_BYTE_WIDTH 4
`define BLOCK_0_REGISTER_3_BYTE_SIZE 4
`define BLOCK_0_REGISTER_3_BYTE_OFFSET 8'h08
`define BLOCK_0_REGISTER_4_BIT_FIELD_0_BIT_WIDTH 4
`define BLOCK_0_REGISTER_4_BIT_FIELD_0_BIT_MASK 4'hf
`define BLOCK_0_REGISTER_4_BIT_FIELD_0_BIT_OFFSET 0
`define BLOCK_0_REGISTER_4_BIT_FIELD_1_BIT_WIDTH 4
`define BLOCK_0_REGISTER_4_BIT_FIELD_1_BIT_MASK 4'hf
`define BLOCK_0_REGISTER_4_BIT_FIELD_1_BIT_OFFSET 8
`define BLOCK_0_REGISTER_4_BIT_FIELD_2_BIT_WIDTH 4
`define BLOCK_0_REGISTER_4_BIT_FIELD_2_BIT_MASK 4'hf
`define BLOCK_0_REGISTER_4_BIT_FIELD_2_BIT_OFFSET 12
`define BLOCK_0_REGISTER_4_BIT_FIELD_3_BIT_WIDTH 4
`define BLOCK_0_REGISTER_4_BIT_FIELD_3_BIT_MASK 4'hf
`define BLOCK_0_REGISTER_4_BIT_FIELD_3_BIT_OFFSET 16
`define BLOCK_0_REGISTER_4_BYTE_WIDTH 4
`define BLOCK_0_REGISTER_4_BYTE_SIZE 4
`define BLOCK_0_REGISTER_4_BYTE_OFFSET 8'h0c
`define BLOCK_0_REGISTER_5_BIT_FIELD_0_BIT_WIDTH 2
`define BLOCK_0_REGISTER_5_BIT_FIELD_0_BIT_MASK 2'h3
`define BLOCK_0_REGISTER_5_BIT_FIELD_0_BIT_OFFSET 0
`define BLOCK_0_REGISTER_5_BIT_FIELD_1_BIT_WIDTH 2
`define BLOCK_0_REGISTER_5_BIT_FIELD_1_BIT_MASK 2'h3
`define BLOCK_0_REGISTER_5_BIT_FIELD_1_BIT_OFFSET 2
`define BLOCK_0_REGISTER_5_BIT_FIELD_2_BIT_WIDTH 2
`define BLOCK_0_REGISTER_5_BIT_FIELD_2_BIT_MASK 2'h3
`define BLOCK_0_REGISTER_5_BIT_FIELD_2_BIT_OFFSET 4
`define BLOCK_0_REGISTER_5_BIT_FIELD_3_BIT_WIDTH 2
`define BLOCK_0_REGISTER_5_BIT_FIELD_3_BIT_MASK 2'h3
`define BLOCK_0_REGISTER_5_BIT_FIELD_3_BIT_OFFSET 6
`define BLOCK_0_REGISTER_5_BIT_FIELD_4_BIT_WIDTH 2
`define BLOCK_0_REGISTER_5_BIT_FIELD_4_BIT_MASK 2'h3
`define BLOCK_0_REGISTER_5_BIT_FIELD_4_BIT_OFFSET 8
`define BLOCK_0_REGISTER_5_BIT_FIELD_5_BIT_WIDTH 2
`define BLOCK_0_REGISTER_5_BIT_FIELD_5_BIT_MASK 2'h3
`define BLOCK_0_REGISTER_5_BIT_FIELD_5_BIT_OFFSET 10
`define BLOCK_0_REGISTER_5_BIT_FIELD_6_BIT_WIDTH 2
`define BLOCK_0_REGISTER_5_BIT_FIELD_6_BIT_MASK 2'h3
`define BLOCK_0_REGISTER_5_BIT_FIELD_6_BIT_OFFSET 12
`define BLOCK_0_REGISTER_5_BIT_FIELD_7_BIT_WIDTH 2
`define BLOCK_0_REGISTER_5_BIT_FIELD_7_BIT_MASK 2'h3
`define BLOCK_0_REGISTER_5_BIT_FIELD_7_BIT_OFFSET 16
`define BLOCK_0_REGISTER_5_BIT_FIELD_8_BIT_WIDTH 2
`define BLOCK_0_REGISTER_5_BIT_FIELD_8_BIT_MASK 2'h3
`define BLOCK_0_REGISTER_5_BIT_FIELD_8_BIT_OFFSET 18
`define BLOCK_0_REGISTER_5_BIT_FIELD_9_BIT_WIDTH 2
`define BLOCK_0_REGISTER_5_BIT_FIELD_9_BIT_MASK 2'h3
`define BLOCK_0_REGISTER_5_BIT_FIELD_9_BIT_OFFSET 20
`define BLOCK_0_REGISTER_5_BYTE_WIDTH 4
`define BLOCK_0_REGISTER_5_BYTE_SIZE 4
`define BLOCK_0_REGISTER_5_BYTE_OFFSET 8'h10
`define BLOCK_0_REGISTER_6_BIT_FIELD_0_BIT_WIDTH 4
`define BLOCK_0_REGISTER_6_BIT_FIELD_0_BIT_MASK 4'hf
`define BLOCK_0_REGISTER_6_BIT_FIELD_0_BIT_OFFSET 0
`define BLOCK_0_REGISTER_6_BIT_FIELD_1_BIT_WIDTH 4
`define BLOCK_0_REGISTER_6_BIT_FIELD_1_BIT_MASK 4'hf
`define BLOCK_0_REGISTER_6_BIT_FIELD_1_BIT_OFFSET 4
`define BLOCK_0_REGISTER_6_BIT_FIELD_2_BIT_WIDTH 4
`define BLOCK_0_REGISTER_6_BIT_FIELD_2_BIT_MASK 4'hf
`define BLOCK_0_REGISTER_6_BIT_FIELD_2_BIT_OFFSET 8
`define BLOCK_0_REGISTER_6_BIT_FIELD_3_BIT_WIDTH 4
`define BLOCK_0_REGISTER_6_BIT_FIELD_3_BIT_MASK 4'hf
`define BLOCK_0_REGISTER_6_BIT_FIELD_3_BIT_OFFSET 12
`define BLOCK_0_REGISTER_6_BIT_FIELD_4_BIT_WIDTH 4
`define BLOCK_0_REGISTER_6_BIT_FIELD_4_BIT_MASK 4'hf
`define BLOCK_0_REGISTER_6_BIT_FIELD_4_BIT_OFFSET 16
`define BLOCK_0_REGISTER_6_BIT_FIELD_5_BIT_WIDTH 4
`define BLOCK_0_REGISTER_6_BIT_FIELD_5_BIT_MASK 4'hf
`define BLOCK_0_REGISTER_6_BIT_FIELD_5_BIT_OFFSET 20
`define BLOCK_0_REGISTER_6_BIT_FIELD_6_BIT_WIDTH 4
`define BLOCK_0_REGISTER_6_BIT_FIELD_6_BIT_MASK 4'hf
`define BLOCK_0_REGISTER_6_BIT_FIELD_6_BIT_OFFSET 24
`define BLOCK_0_REGISTER_6_BIT_FIELD_7_BIT_WIDTH 4
`define BLOCK_0_REGISTER_6_BIT_FIELD_7_BIT_MASK 4'hf
`define BLOCK_0_REGISTER_6_BIT_FIELD_7_BIT_OFFSET 28
`define BLOCK_0_REGISTER_6_BIT_FIELD_8_BIT_WIDTH 4
`define BLOCK_0_REGISTER_6_BIT_FIELD_8_BIT_MASK 4'hf
`define BLOCK_0_REGISTER_6_BIT_FIELD_8_BIT_OFFSET 32
`define BLOCK_0_REGISTER_6_BIT_FIELD_9_BIT_WIDTH 4
`define BLOCK_0_REGISTER_6_BIT_FIELD_9_BIT_MASK 4'hf
`define BLOCK_0_REGISTER_6_BIT_FIELD_9_BIT_OFFSET 36
`define BLOCK_0_REGISTER_6_BYTE_WIDTH 8
`define BLOCK_0_REGISTER_6_BYTE_SIZE 8
`define BLOCK_0_REGISTER_6_BYTE_OFFSET 8'h14
`define BLOCK_0_REGISTER_7_BIT_FIELD_0_BIT_WIDTH 4
`define BLOCK_0_REGISTER_7_BIT_FIELD_0_BIT_MASK 4'hf
`define BLOCK_0_REGISTER_7_BIT_FIELD_0_BIT_OFFSET 0
`define BLOCK_0_REGISTER_7_BIT_FIELD_1_BIT_WIDTH 4
`define BLOCK_0_REGISTER_7_BIT_FIELD_1_BIT_MASK 4'hf
`define BLOCK_0_REGISTER_7_BIT_FIELD_1_BIT_OFFSET 8
`define BLOCK_0_REGISTER_7_BIT_FIELD_2_BIT_WIDTH 4
`define BLOCK_0_REGISTER_7_BIT_FIELD_2_BIT_MASK 4'hf
`define BLOCK_0_REGISTER_7_BIT_FIELD_2_BIT_OFFSET 16
`define BLOCK_0_REGISTER_7_BIT_FIELD_3_BIT_WIDTH 4
`define BLOCK_0_REGISTER_7_BIT_FIELD_3_BIT_MASK 4'hf
`define BLOCK_0_REGISTER_7_BIT_FIELD_3_BIT_OFFSET 24
`define BLOCK_0_REGISTER_7_BYTE_WIDTH 4
`define BLOCK_0_REGISTER_7_BYTE_SIZE 4
`define BLOCK_0_REGISTER_7_BYTE_OFFSET 8'h1c
`define BLOCK_0_REGISTER_8_BIT_FIELD_0_BIT_WIDTH 4
`define BLOCK_0_REGISTER_8_BIT_FIELD_0_BIT_MASK 4'hf
`define BLOCK_0_REGISTER_8_BIT_FIELD_0_BIT_OFFSET 0
`define BLOCK_0_REGISTER_8_BIT_FIELD_1_BIT_WIDTH 4
`define BLOCK_0_REGISTER_8_BIT_FIELD_1_BIT_MASK 4'hf
`define BLOCK_0_REGISTER_8_BIT_FIELD_1_BIT_OFFSET 8
`define BLOCK_0_REGISTER_8_BIT_FIELD_2_BIT_WIDTH 4
`define BLOCK_0_REGISTER_8_BIT_FIELD_2_BIT_MASK 4'hf
`define BLOCK_0_REGISTER_8_BIT_FIELD_2_BIT_OFFSET 16
`define BLOCK_0_REGISTER_8_BIT_FIELD_3_BIT_WIDTH 4
`define BLOCK_0_REGISTER_8_BIT_FIELD_3_BIT_MASK 4'hf
`define BLOCK_0_REGISTER_8_BIT_FIELD_3_BIT_OFFSET 24
`define BLOCK_0_REGISTER_8_BIT_FIELD_4_BIT_WIDTH 4
`define BLOCK_0_REGISTER_8_BIT_FIELD_4_BIT_MASK 4'hf
`define BLOCK_0_REGISTER_8_BIT_FIELD_4_BIT_OFFSET 32
`define BLOCK_0_REGISTER_8_BIT_FIELD_5_BIT_WIDTH 4
`define BLOCK_0_REGISTER_8_BIT_FIELD_5_BIT_MASK 4'hf
`define BLOCK_0_REGISTER_8_BIT_FIELD_5_BIT_OFFSET 40
`define BLOCK_0_REGISTER_8_BYTE_WIDTH 8
`define BLOCK_0_REGISTER_8_BYTE_SIZE 8
`define BLOCK_0_REGISTER_8_BYTE_OFFSET 8'h20
`define BLOCK_0_REGISTER_9_BIT_FIELD_0_BIT_WIDTH 2
`define BLOCK_0_REGISTER_9_BIT_FIELD_0_BIT_MASK 2'h3
`define BLOCK_0_REGISTER_9_BIT_FIELD_0_BIT_OFFSET 0
`define BLOCK_0_REGISTER_9_BIT_FIELD_1_BIT_WIDTH 2
`define BLOCK_0_REGISTER_9_BIT_FIELD_1_BIT_MASK 2'h3
`define BLOCK_0_REGISTER_9_BIT_FIELD_1_BIT_OFFSET 2
`define BLOCK_0_REGISTER_9_BIT_FIELD_2_BIT_WIDTH 2
`define BLOCK_0_REGISTER_9_BIT_FIELD_2_BIT_MASK 2'h3
`define BLOCK_0_REGISTER_9_BIT_FIELD_2_BIT_OFFSET 4
`define BLOCK_0_REGISTER_9_BIT_FIELD_3_BIT_WIDTH 2
`define BLOCK_0_REGISTER_9_BIT_FIELD_3_BIT_MASK 2'h3
`define BLOCK_0_REGISTER_9_BIT_FIELD_3_BIT_OFFSET 6
`define BLOCK_0_REGISTER_9_BIT_FIELD_4_BIT_WIDTH 2
`define BLOCK_0_REGISTER_9_BIT_FIELD_4_BIT_MASK 2'h3
`define BLOCK_0_REGISTER_9_BIT_FIELD_4_BIT_OFFSET 8
`define BLOCK_0_REGISTER_9_BIT_FIELD_5_BIT_WIDTH 2
`define BLOCK_0_REGISTER_9_BIT_FIELD_5_BIT_MASK 2'h3
`define BLOCK_0_REGISTER_9_BIT_FIELD_5_BIT_OFFSET 10
`define BLOCK_0_REGISTER_9_BYTE_WIDTH 4
`define BLOCK_0_REGISTER_9_BYTE_SIZE 4
`define BLOCK_0_REGISTER_9_BYTE_OFFSET 8'h28
`define BLOCK_0_REGISTER_10_BIT_FIELD_0_BIT_WIDTH 2
`define BLOCK_0_REGISTER_10_BIT_FIELD_0_BIT_MASK 2'h3
`define BLOCK_0_REGISTER_10_BIT_FIELD_0_BIT_OFFSET_0 0
`define BLOCK_0_REGISTER_10_BIT_FIELD_0_BIT_OFFSET_1 8
`define BLOCK_0_REGISTER_10_BIT_FIELD_0_BIT_OFFSET_2 16
`define BLOCK_0_REGISTER_10_BIT_FIELD_0_BIT_OFFSET_3 24
`define BLOCK_0_REGISTER_10_BIT_FIELD_1_BIT_WIDTH 2
`define BLOCK_0_REGISTER_10_BIT_FIELD_1_BIT_MASK 2'h3
`define BLOCK_0_REGISTER_10_BIT_FIELD_1_BIT_OFFSET_0 2
`define BLOCK_0_REGISTER_10_BIT_FIELD_1_BIT_OFFSET_1 10
`define BLOCK_0_REGISTER_10_BIT_FIELD_1_BIT_OFFSET_2 18
`define BLOCK_0_REGISTER_10_BIT_FIELD_1_BIT_OFFSET_3 26
`define BLOCK_0_REGISTER_10_BIT_FIELD_2_BIT_WIDTH 2
`define BLOCK_0_REGISTER_10_BIT_FIELD_2_BIT_MASK 2'h3
`define BLOCK_0_REGISTER_10_BIT_FIELD_2_BIT_OFFSET_0 4
`define BLOCK_0_REGISTER_10_BIT_FIELD_2_BIT_OFFSET_1 12
`define BLOCK_0_REGISTER_10_BIT_FIELD_2_BIT_OFFSET_2 20
`define BLOCK_0_REGISTER_10_BIT_FIELD_2_BIT_OFFSET_3 28
`define BLOCK_0_REGISTER_10_BYTE_WIDTH 4
`define BLOCK_0_REGISTER_10_BYTE_SIZE 32
`define BLOCK_0_REGISTER_10_ARRAY_DIMENSION 1
`define BLOCK_0_REGISTER_10_ARRAY_SIZE_0 4
`define BLOCK_0_REGISTER_10_BYTE_OFFSET_0 8'h30
`define BLOCK_0_REGISTER_10_BYTE_OFFSET_1 8'h38
`define BLOCK_0_REGISTER_10_BYTE_OFFSET_2 8'h40
`define BLOCK_0_REGISTER_10_BYTE_OFFSET_3 8'h48
`define BLOCK_0_REGISTER_11_BIT_FIELD_0_BIT_WIDTH 8
`define BLOCK_0_REGISTER_11_BIT_FIELD_0_BIT_MASK 8'hff
`define BLOCK_0_REGISTER_11_BIT_FIELD_0_BIT_OFFSET_0 0
`define BLOCK_0_REGISTER_11_BIT_FIELD_0_BIT_OFFSET_1 16
`define BLOCK_0_REGISTER_11_BIT_FIELD_0_BIT_OFFSET_2 32
`define BLOCK_0_REGISTER_11_BIT_FIELD_0_BIT_OFFSET_3 48
`define BLOCK_0_REGISTER_11_BIT_FIELD_1_BIT_WIDTH 8
`define BLOCK_0_REGISTER_11_BIT_FIELD_1_BIT_MASK 8'hff
`define BLOCK_0_REGISTER_11_BIT_FIELD_1_BIT_OFFSET_0 8
`define BLOCK_0_REGISTER_11_BIT_FIELD_1_BIT_OFFSET_1 24
`define BLOCK_0_REGISTER_11_BIT_FIELD_1_BIT_OFFSET_2 40
`define BLOCK_0_REGISTER_11_BIT_FIELD_1_BIT_OFFSET_3 56
`define BLOCK_0_REGISTER_11_BYTE_WIDTH 8
`define BLOCK_0_REGISTER_11_BYTE_SIZE 8
`define BLOCK_0_REGISTER_11_ARRAY_DIMENSION 2
`define BLOCK_0_REGISTER_11_ARRAY_SIZE_0 2
`define BLOCK_0_REGISTER_11_ARRAY_SIZE_1 4
`define BLOCK_0_REGISTER_11_BYTE_OFFSET_0_0 8'h50
`define BLOCK_0_REGISTER_11_BYTE_OFFSET_0_1 8'h50
`define BLOCK_0_REGISTER_11_BYTE_OFFSET_0_2 8'h50
`define BLOCK_0_REGISTER_11_BYTE_OFFSET_0_3 8'h50
`define BLOCK_0_REGISTER_11_BYTE_OFFSET_1_0 8'h50
`define BLOCK_0_REGISTER_11_BYTE_OFFSET_1_1 8'h50
`define BLOCK_0_REGISTER_11_BYTE_OFFSET_1_2 8'h50
`define BLOCK_0_REGISTER_11_BYTE_OFFSET_1_3 8'h50
`define BLOCK_0_REGISTER_12_BIT_FIELD_0_BIT_WIDTH 1
`define BLOCK_0_REGISTER_12_BIT_FIELD_0_BIT_MASK 1'h1
`define BLOCK_0_REGISTER_12_BIT_FIELD_0_BIT_OFFSET 0
`define BLOCK_0_REGISTER_12_BIT_FIELD_1_BIT_WIDTH 1
`define BLOCK_0_REGISTER_12_BIT_FIELD_1_BIT_MASK 1'h1
`define BLOCK_0_REGISTER_12_BIT_FIELD_1_BIT_OFFSET 32
`define BLOCK_0_REGISTER_12_BYTE_WIDTH 8
`define BLOCK_0_REGISTER_12_BYTE_SIZE 8
`define BLOCK_0_REGISTER_12_BYTE_OFFSET 8'h50
`define BLOCK_0_REGISTER_13_BIT_FIELD_0_BIT_WIDTH 2
`define BLOCK_0_REGISTER_13_BIT_FIELD_0_BIT_MASK 2'h3
`define BLOCK_0_REGISTER_13_BIT_FIELD_0_BIT_OFFSET 0
`define BLOCK_0_REGISTER_13_BIT_FIELD_1_BIT_WIDTH 2
`define BLOCK_0_REGISTER_13_BIT_FIELD_1_BIT_MASK 2'h3
`define BLOCK_0_REGISTER_13_BIT_FIELD_1_BIT_OFFSET 2
`define BLOCK_0_REGISTER_13_BIT_FIELD_2_BIT_WIDTH 2
`define BLOCK_0_REGISTER_13_BIT_FIELD_2_BIT_MASK 2'h3
`define BLOCK_0_REGISTER_13_BIT_FIELD_2_BIT_OFFSET 4
`define BLOCK_0_REGISTER_13_BIT_FIELD_3_BIT_WIDTH 2
`define BLOCK_0_REGISTER_13_BIT_FIELD_3_BIT_MASK 2'h3
`define BLOCK_0_REGISTER_13_BIT_FIELD_3_BIT_OFFSET 6
`define BLOCK_0_REGISTER_13_BIT_FIELD_4_BIT_WIDTH 2
`define BLOCK_0_REGISTER_13_BIT_FIELD_4_BIT_MASK 2'h3
`define BLOCK_0_REGISTER_13_BIT_FIELD_4_BIT_OFFSET 8
`define BLOCK_0_REGISTER_13_BIT_FIELD_5_BIT_WIDTH 2
`define BLOCK_0_REGISTER_13_BIT_FIELD_5_BIT_MASK 2'h3
`define BLOCK_0_REGISTER_13_BIT_FIELD_5_BIT_OFFSET 10
`define BLOCK_0_REGISTER_13_BIT_FIELD_6_BIT_WIDTH 2
`define BLOCK_0_REGISTER_13_BIT_FIELD_6_BIT_MASK 2'h3
`define BLOCK_0_REGISTER_13_BIT_FIELD_6_BIT_OFFSET 12
`define BLOCK_0_REGISTER_13_BIT_FIELD_7_BIT_WIDTH 2
`define BLOCK_0_REGISTER_13_BIT_FIELD_7_BIT_MASK 2'h3
`define BLOCK_0_REGISTER_13_BIT_FIELD_7_BIT_OFFSET 14
`define BLOCK_0_REGISTER_13_BIT_FIELD_8_BIT_WIDTH 2
`define BLOCK_0_REGISTER_13_BIT_FIELD_8_BIT_MASK 2'h3
`define BLOCK_0_REGISTER_13_BIT_FIELD_8_BIT_OFFSET 16
`define BLOCK_0_REGISTER_13_BYTE_WIDTH 4
`define BLOCK_0_REGISTER_13_BYTE_SIZE 4
`define BLOCK_0_REGISTER_13_BYTE_OFFSET 8'h60
`define BLOCK_0_REGISTER_14_BIT_FIELD_0_BIT_WIDTH 1
`define BLOCK_0_REGISTER_14_BIT_FIELD_0_BIT_MASK 1'h1
`define BLOCK_0_REGISTER_14_BIT_FIELD_0_BIT_OFFSET 0
`define BLOCK_0_REGISTER_14_BYTE_WIDTH 4
`define BLOCK_0_REGISTER_14_BYTE_SIZE 4
`define BLOCK_0_REGISTER_14_BYTE_OFFSET 8'h70
`define BLOCK_0_REGISTER_15_BIT_FIELD_0_BIT_WIDTH 1
`define BLOCK_0_REGISTER_15_BIT_FIELD_0_BIT_MASK 1'h1
`define BLOCK_0_REGISTER_15_BIT_FIELD_0_BIT_OFFSET 0
`define BLOCK_0_REGISTER_15_BYTE_WIDTH 4
`define BLOCK_0_REGISTER_15_BYTE_SIZE 4
`define BLOCK_0_REGISTER_15_BYTE_OFFSET 8'h74
`define BLOCK_0_REGISTER_17_BYTE_WIDTH 4
`define BLOCK_0_REGISTER_17_BYTE_SIZE 128
`define BLOCK_0_REGISTER_17_BYTE_OFFSET 8'h80
`endif
