package uart_csr_rtl_pkg;
  localparam int RBR_BYTE_WIDTH = 4;
  localparam int RBR_BYTE_SIZE = 4;
  localparam bit [4:0] RBR_BYTE_OFFSET = 5'h00;
  localparam int RBR_BIT_WIDTH = 8;
  localparam bit [7:0] RBR_BIT_MASK = 8'hff;
  localparam int RBR_BIT_OFFSET = 0;
  localparam int THR_BYTE_WIDTH = 4;
  localparam int THR_BYTE_SIZE = 4;
  localparam bit [4:0] THR_BYTE_OFFSET = 5'h00;
  localparam int THR_BIT_WIDTH = 8;
  localparam bit [7:0] THR_BIT_MASK = 8'hff;
  localparam int THR_BIT_OFFSET = 0;
  localparam int IER_BYTE_WIDTH = 4;
  localparam int IER_BYTE_SIZE = 4;
  localparam bit [4:0] IER_BYTE_OFFSET = 5'h04;
  localparam int IER_ERBFI_BIT_WIDTH = 1;
  localparam bit IER_ERBFI_BIT_MASK = 1'h1;
  localparam int IER_ERBFI_BIT_OFFSET = 0;
  localparam int IER_ETBEI_BIT_WIDTH = 1;
  localparam bit IER_ETBEI_BIT_MASK = 1'h1;
  localparam int IER_ETBEI_BIT_OFFSET = 1;
  localparam int IER_ELSI_BIT_WIDTH = 1;
  localparam bit IER_ELSI_BIT_MASK = 1'h1;
  localparam int IER_ELSI_BIT_OFFSET = 2;
  localparam int IER_EDSSI_BIT_WIDTH = 1;
  localparam bit IER_EDSSI_BIT_MASK = 1'h1;
  localparam int IER_EDSSI_BIT_OFFSET = 3;
  localparam int IIR_BYTE_WIDTH = 4;
  localparam int IIR_BYTE_SIZE = 4;
  localparam bit [4:0] IIR_BYTE_OFFSET = 5'h08;
  localparam int IIR_INTPEND_BIT_WIDTH = 1;
  localparam bit IIR_INTPEND_BIT_MASK = 1'h1;
  localparam int IIR_INTPEND_BIT_OFFSET = 0;
  localparam int IIR_INTID2_BIT_WIDTH = 3;
  localparam bit [2:0] IIR_INTID2_BIT_MASK = 3'h7;
  localparam int IIR_INTID2_BIT_OFFSET = 1;
  localparam int FCR_BYTE_WIDTH = 4;
  localparam int FCR_BYTE_SIZE = 4;
  localparam bit [4:0] FCR_BYTE_OFFSET = 5'h08;
  localparam int FCR_FIFOEN_BIT_WIDTH = 1;
  localparam bit FCR_FIFOEN_BIT_MASK = 1'h1;
  localparam int FCR_FIFOEN_BIT_OFFSET = 0;
  localparam int FCR_RCVR_FIFO_RESET_BIT_WIDTH = 1;
  localparam bit FCR_RCVR_FIFO_RESET_BIT_MASK = 1'h1;
  localparam int FCR_RCVR_FIFO_RESET_BIT_OFFSET = 1;
  localparam int FCR_XMIT_FIFO_RESET_BIT_WIDTH = 1;
  localparam bit FCR_XMIT_FIFO_RESET_BIT_MASK = 1'h1;
  localparam int FCR_XMIT_FIFO_RESET_BIT_OFFSET = 2;
  localparam int FCR_DMA_MODE_SELECT_BIT_WIDTH = 1;
  localparam bit FCR_DMA_MODE_SELECT_BIT_MASK = 1'h1;
  localparam int FCR_DMA_MODE_SELECT_BIT_OFFSET = 3;
  localparam int FCR_RCVR_FIFO_TRIGGER_LEVEL_BIT_WIDTH = 2;
  localparam bit [1:0] FCR_RCVR_FIFO_TRIGGER_LEVEL_BIT_MASK = 2'h3;
  localparam int FCR_RCVR_FIFO_TRIGGER_LEVEL_BIT_OFFSET = 6;
  localparam int LCR_BYTE_WIDTH = 4;
  localparam int LCR_BYTE_SIZE = 4;
  localparam bit [4:0] LCR_BYTE_OFFSET = 5'h0c;
  localparam int LCR_WLS_BIT_WIDTH = 2;
  localparam bit [1:0] LCR_WLS_BIT_MASK = 2'h3;
  localparam int LCR_WLS_BIT_OFFSET = 0;
  localparam int LCR_STB_BIT_WIDTH = 1;
  localparam bit LCR_STB_BIT_MASK = 1'h1;
  localparam int LCR_STB_BIT_OFFSET = 2;
  localparam int LCR_PEN_BIT_WIDTH = 1;
  localparam bit LCR_PEN_BIT_MASK = 1'h1;
  localparam int LCR_PEN_BIT_OFFSET = 3;
  localparam int LCR_EPS_BIT_WIDTH = 1;
  localparam bit LCR_EPS_BIT_MASK = 1'h1;
  localparam int LCR_EPS_BIT_OFFSET = 4;
  localparam int LCR_STICK_PARITY_BIT_WIDTH = 1;
  localparam bit LCR_STICK_PARITY_BIT_MASK = 1'h1;
  localparam int LCR_STICK_PARITY_BIT_OFFSET = 5;
  localparam int LCR_SET_BREAK_BIT_WIDTH = 1;
  localparam bit LCR_SET_BREAK_BIT_MASK = 1'h1;
  localparam int LCR_SET_BREAK_BIT_OFFSET = 6;
  localparam int LCR_DLAB_BIT_WIDTH = 1;
  localparam bit LCR_DLAB_BIT_MASK = 1'h1;
  localparam int LCR_DLAB_BIT_OFFSET = 7;
  localparam int MRC_BYTE_WIDTH = 4;
  localparam int MRC_BYTE_SIZE = 4;
  localparam bit [4:0] MRC_BYTE_OFFSET = 5'h10;
  localparam int MRC_DTR_BIT_WIDTH = 1;
  localparam bit MRC_DTR_BIT_MASK = 1'h1;
  localparam int MRC_DTR_BIT_OFFSET = 0;
  localparam int MRC_RTS_BIT_WIDTH = 1;
  localparam bit MRC_RTS_BIT_MASK = 1'h1;
  localparam int MRC_RTS_BIT_OFFSET = 1;
  localparam int MRC_OUT1_BIT_WIDTH = 1;
  localparam bit MRC_OUT1_BIT_MASK = 1'h1;
  localparam int MRC_OUT1_BIT_OFFSET = 2;
  localparam int MRC_OUT2_BIT_WIDTH = 1;
  localparam bit MRC_OUT2_BIT_MASK = 1'h1;
  localparam int MRC_OUT2_BIT_OFFSET = 3;
  localparam int MRC_LOOP_BACK_BIT_WIDTH = 1;
  localparam bit MRC_LOOP_BACK_BIT_MASK = 1'h1;
  localparam int MRC_LOOP_BACK_BIT_OFFSET = 4;
  localparam int LSR_BYTE_WIDTH = 4;
  localparam int LSR_BYTE_SIZE = 4;
  localparam bit [4:0] LSR_BYTE_OFFSET = 5'h14;
  localparam int LSR_DR_BIT_WIDTH = 1;
  localparam bit LSR_DR_BIT_MASK = 1'h1;
  localparam int LSR_DR_BIT_OFFSET = 0;
  localparam int LSR_OE_BIT_WIDTH = 1;
  localparam bit LSR_OE_BIT_MASK = 1'h1;
  localparam int LSR_OE_BIT_OFFSET = 1;
  localparam int LSR_PE_BIT_WIDTH = 1;
  localparam bit LSR_PE_BIT_MASK = 1'h1;
  localparam int LSR_PE_BIT_OFFSET = 2;
  localparam int LSR_FE_BIT_WIDTH = 1;
  localparam bit LSR_FE_BIT_MASK = 1'h1;
  localparam int LSR_FE_BIT_OFFSET = 3;
  localparam int LSR_BI_BIT_WIDTH = 1;
  localparam bit LSR_BI_BIT_MASK = 1'h1;
  localparam int LSR_BI_BIT_OFFSET = 4;
  localparam int LSR_THRE_BIT_WIDTH = 1;
  localparam bit LSR_THRE_BIT_MASK = 1'h1;
  localparam int LSR_THRE_BIT_OFFSET = 5;
  localparam int LSR_TEMT_BIT_WIDTH = 1;
  localparam bit LSR_TEMT_BIT_MASK = 1'h1;
  localparam int LSR_TEMT_BIT_OFFSET = 6;
  localparam int LSR_ERROR_IN_RCVR_FIFO_BIT_WIDTH = 1;
  localparam bit LSR_ERROR_IN_RCVR_FIFO_BIT_MASK = 1'h1;
  localparam int LSR_ERROR_IN_RCVR_FIFO_BIT_OFFSET = 7;
  localparam int MSR_BYTE_WIDTH = 4;
  localparam int MSR_BYTE_SIZE = 4;
  localparam bit [4:0] MSR_BYTE_OFFSET = 5'h18;
  localparam int MSR_DCTS_BIT_WIDTH = 1;
  localparam bit MSR_DCTS_BIT_MASK = 1'h1;
  localparam int MSR_DCTS_BIT_OFFSET = 0;
  localparam int MSR_DDSR_BIT_WIDTH = 1;
  localparam bit MSR_DDSR_BIT_MASK = 1'h1;
  localparam int MSR_DDSR_BIT_OFFSET = 1;
  localparam int MSR_TERI_BIT_WIDTH = 1;
  localparam bit MSR_TERI_BIT_MASK = 1'h1;
  localparam int MSR_TERI_BIT_OFFSET = 2;
  localparam int MSR_DDCD_BIT_WIDTH = 1;
  localparam bit MSR_DDCD_BIT_MASK = 1'h1;
  localparam int MSR_DDCD_BIT_OFFSET = 3;
  localparam int MSR_CTS_BIT_WIDTH = 1;
  localparam bit MSR_CTS_BIT_MASK = 1'h1;
  localparam int MSR_CTS_BIT_OFFSET = 4;
  localparam int MSR_DSR_BIT_WIDTH = 1;
  localparam bit MSR_DSR_BIT_MASK = 1'h1;
  localparam int MSR_DSR_BIT_OFFSET = 5;
  localparam int MSR_RI_BIT_WIDTH = 1;
  localparam bit MSR_RI_BIT_MASK = 1'h1;
  localparam int MSR_RI_BIT_OFFSET = 6;
  localparam int MSR_DCD_BIT_WIDTH = 1;
  localparam bit MSR_DCD_BIT_MASK = 1'h1;
  localparam int MSR_DCD_BIT_OFFSET = 7;
  localparam int SCRATCH_BYTE_WIDTH = 4;
  localparam int SCRATCH_BYTE_SIZE = 4;
  localparam bit [4:0] SCRATCH_BYTE_OFFSET = 5'h1c;
  localparam int SCRATCH_BIT_WIDTH = 8;
  localparam bit [7:0] SCRATCH_BIT_MASK = 8'hff;
  localparam int SCRATCH_BIT_OFFSET = 0;
  localparam int DLL_BYTE_WIDTH = 4;
  localparam int DLL_BYTE_SIZE = 4;
  localparam bit [4:0] DLL_BYTE_OFFSET = 5'h00;
  localparam int DLL_BIT_WIDTH = 8;
  localparam bit [7:0] DLL_BIT_MASK = 8'hff;
  localparam int DLL_BIT_OFFSET = 0;
  localparam int DLM_BYTE_WIDTH = 4;
  localparam int DLM_BYTE_SIZE = 4;
  localparam bit [4:0] DLM_BYTE_OFFSET = 5'h04;
  localparam int DLM_BIT_WIDTH = 8;
  localparam bit [7:0] DLM_BIT_MASK = 8'hff;
  localparam int DLM_BIT_OFFSET = 0;
endpackage
