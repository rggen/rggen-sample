`ifndef BLOCK_1_VH
`define BLOCK_1_VH
`define BLOCK_1_REGISTER_FILE_0_REGISTER_0_BIT_FIELD_0_BIT_WIDTH 8
`define BLOCK_1_REGISTER_FILE_0_REGISTER_0_BIT_FIELD_0_BIT_MASK 8'hff
`define BLOCK_1_REGISTER_FILE_0_REGISTER_0_BIT_FIELD_0_BIT_OFFSET 0
`define BLOCK_1_REGISTER_FILE_0_REGISTER_0_BYTE_WIDTH 4
`define BLOCK_1_REGISTER_FILE_0_REGISTER_0_BYTE_SIZE 4
`define BLOCK_1_REGISTER_FILE_0_REGISTER_0_BYTE_OFFSET 7'h00
`define BLOCK_1_REGISTER_FILE_0_REGISTER_1_BIT_FIELD_0_BIT_WIDTH 8
`define BLOCK_1_REGISTER_FILE_0_REGISTER_1_BIT_FIELD_0_BIT_MASK 8'hff
`define BLOCK_1_REGISTER_FILE_0_REGISTER_1_BIT_FIELD_0_BIT_OFFSET 0
`define BLOCK_1_REGISTER_FILE_0_REGISTER_1_BYTE_WIDTH 4
`define BLOCK_1_REGISTER_FILE_0_REGISTER_1_BYTE_SIZE 4
`define BLOCK_1_REGISTER_FILE_0_REGISTER_1_BYTE_OFFSET 7'h04
`define BLOCK_1_REGISTER_FILE_1_REGISTER_0_BIT_FIELD_0_BIT_WIDTH 8
`define BLOCK_1_REGISTER_FILE_1_REGISTER_0_BIT_FIELD_0_BIT_MASK 8'hff
`define BLOCK_1_REGISTER_FILE_1_REGISTER_0_BIT_FIELD_0_BIT_OFFSET 0
`define BLOCK_1_REGISTER_FILE_1_REGISTER_0_BYTE_WIDTH 4
`define BLOCK_1_REGISTER_FILE_1_REGISTER_0_BYTE_SIZE 4
`define BLOCK_1_REGISTER_FILE_1_REGISTER_0_ARRAY_DIMENSION 1
`define BLOCK_1_REGISTER_FILE_1_REGISTER_0_ARRAY_SIZE_0 2
`define BLOCK_1_REGISTER_FILE_1_REGISTER_0_BYTE_OFFSET_0 7'h10
`define BLOCK_1_REGISTER_FILE_1_REGISTER_0_BYTE_OFFSET_1 7'h10
`define BLOCK_1_REGISTER_FILE_1_REGISTER_1_BIT_FIELD_0_BIT_WIDTH 8
`define BLOCK_1_REGISTER_FILE_1_REGISTER_1_BIT_FIELD_0_BIT_MASK 8'hff
`define BLOCK_1_REGISTER_FILE_1_REGISTER_1_BIT_FIELD_0_BIT_OFFSET 0
`define BLOCK_1_REGISTER_FILE_1_REGISTER_1_BYTE_WIDTH 4
`define BLOCK_1_REGISTER_FILE_1_REGISTER_1_BYTE_SIZE 4
`define BLOCK_1_REGISTER_FILE_1_REGISTER_1_ARRAY_DIMENSION 1
`define BLOCK_1_REGISTER_FILE_1_REGISTER_1_ARRAY_SIZE_0 2
`define BLOCK_1_REGISTER_FILE_1_REGISTER_1_BYTE_OFFSET_0 7'h10
`define BLOCK_1_REGISTER_FILE_1_REGISTER_1_BYTE_OFFSET_1 7'h10
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_0_BIT_FIELD_0_BIT_WIDTH 4
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_0_BIT_FIELD_0_BIT_MASK 4'hf
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_0_BIT_FIELD_0_BIT_OFFSET_0 0
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_0_BIT_FIELD_0_BIT_OFFSET_1 4
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_0_BIT_FIELD_1_BIT_WIDTH 4
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_0_BIT_FIELD_1_BIT_MASK 4'hf
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_0_BIT_FIELD_1_BIT_OFFSET_0 8
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_0_BIT_FIELD_1_BIT_OFFSET_1 12
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_0_BIT_FIELD_2_BIT_WIDTH 4
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_0_BIT_FIELD_2_BIT_MASK 4'hf
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_0_BIT_FIELD_2_BIT_OFFSET_0 16
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_0_BIT_FIELD_2_BIT_OFFSET_1 20
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_0_BYTE_WIDTH 4
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_0_BYTE_SIZE 48
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_0_ARRAY_DIMENSION 3
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_0_ARRAY_SIZE_0 2
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_0_ARRAY_SIZE_1 2
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_0_ARRAY_SIZE_2 3
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_0_BYTE_OFFSET_0_0_0 7'h20
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_0_BYTE_OFFSET_0_0_1 7'h24
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_0_BYTE_OFFSET_0_0_2 7'h28
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_0_BYTE_OFFSET_0_1_0 7'h2c
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_0_BYTE_OFFSET_0_1_1 7'h30
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_0_BYTE_OFFSET_0_1_2 7'h34
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_0_BYTE_OFFSET_1_0_0 7'h3c
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_0_BYTE_OFFSET_1_0_1 7'h40
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_0_BYTE_OFFSET_1_0_2 7'h44
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_0_BYTE_OFFSET_1_1_0 7'h48
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_0_BYTE_OFFSET_1_1_1 7'h4c
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_0_BYTE_OFFSET_1_1_2 7'h50
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_1_BIT_FIELD_0_BIT_WIDTH 1
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_1_BIT_FIELD_0_BIT_MASK 1'h1
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_1_BIT_FIELD_0_BIT_OFFSET_0 0
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_1_BIT_FIELD_0_BIT_OFFSET_1 1
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_1_BYTE_WIDTH 4
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_1_BYTE_SIZE 8
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_1_ARRAY_DIMENSION 1
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_1_ARRAY_SIZE_0 2
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_1_BYTE_OFFSET_0 7'h38
`define BLOCK_1_REGISTER_FILE_2_REGISTER_FILE_0_REGISTER_1_BYTE_OFFSET_1 7'h54
`endif
