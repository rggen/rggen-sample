package block_0_rtl_pkg;
  localparam int REGISTER_0_BYTE_WIDTH = 4;
  localparam int REGISTER_0_BYTE_SIZE = 4;
  localparam bit [7:0] REGISTER_0_BYTE_OFFSET = 8'h00;
  localparam int REGISTER_0_BIT_FIELD_0_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_0_BIT_FIELD_0_BIT_MASK = 4'hf;
  localparam int REGISTER_0_BIT_FIELD_0_BIT_OFFSET = 0;
  localparam int REGISTER_0_BIT_FIELD_1_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_0_BIT_FIELD_1_BIT_MASK = 4'hf;
  localparam int REGISTER_0_BIT_FIELD_1_BIT_OFFSET = 4;
  localparam int REGISTER_0_BIT_FIELD_2_BIT_WIDTH = 1;
  localparam bit REGISTER_0_BIT_FIELD_2_BIT_MASK = 1'h1;
  localparam int REGISTER_0_BIT_FIELD_2_BIT_OFFSET = 8;
  localparam int REGISTER_0_BIT_FIELD_3_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_0_BIT_FIELD_3_BIT_MASK = 2'h3;
  localparam int REGISTER_0_BIT_FIELD_3_BIT_OFFSET = 9;
  localparam int REGISTER_0_BIT_FIELD_4_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_0_BIT_FIELD_4_BIT_MASK = 2'h3;
  localparam int REGISTER_0_BIT_FIELD_4_BIT_OFFSET = 11;
  localparam int REGISTER_0_BIT_FIELD_5_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_0_BIT_FIELD_5_BIT_MASK = 2'h3;
  localparam int REGISTER_0_BIT_FIELD_5_BIT_OFFSET = 13;
  localparam int REGISTER_0_BIT_FIELD_6_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_0_BIT_FIELD_6_BIT_MASK = 2'h3;
  localparam int REGISTER_0_BIT_FIELD_6_BIT_OFFSET = 15;
  localparam int REGISTER_1_BYTE_WIDTH = 4;
  localparam int REGISTER_1_BYTE_SIZE = 4;
  localparam bit [7:0] REGISTER_1_BYTE_OFFSET = 8'h04;
  localparam int REGISTER_1_BIT_WIDTH = 1;
  localparam bit REGISTER_1_BIT_MASK = 1'h1;
  localparam int REGISTER_1_BIT_OFFSET = 0;
  localparam bit REGISTER_1_FOO = 1'h0;
  localparam bit REGISTER_1_BAR = 1'h1;
  localparam int REGISTER_2_BYTE_WIDTH = 4;
  localparam int REGISTER_2_BYTE_SIZE = 4;
  localparam bit [7:0] REGISTER_2_BYTE_OFFSET = 8'h08;
  localparam int REGISTER_2_BIT_FIELD_0_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_2_BIT_FIELD_0_BIT_MASK = 4'hf;
  localparam int REGISTER_2_BIT_FIELD_0_BIT_OFFSET = 0;
  localparam int REGISTER_2_BIT_FIELD_1_BIT_WIDTH = 8;
  localparam bit [7:0] REGISTER_2_BIT_FIELD_1_BIT_MASK = 8'hff;
  localparam int REGISTER_2_BIT_FIELD_1_BIT_OFFSET = 8;
  localparam int REGISTER_2_BIT_FIELD_2_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_2_BIT_FIELD_2_BIT_MASK = 4'hf;
  localparam int REGISTER_2_BIT_FIELD_2_BIT_OFFSET = 16;
  localparam int REGISTER_2_BIT_FIELD_3_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_2_BIT_FIELD_3_BIT_MASK = 4'hf;
  localparam int REGISTER_2_BIT_FIELD_3_BIT_OFFSET = 20;
  localparam int REGISTER_3_BYTE_WIDTH = 4;
  localparam int REGISTER_3_BYTE_SIZE = 4;
  localparam bit [7:0] REGISTER_3_BYTE_OFFSET = 8'h08;
  localparam int REGISTER_3_BIT_FIELD_0_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_3_BIT_FIELD_0_BIT_MASK = 4'hf;
  localparam int REGISTER_3_BIT_FIELD_0_BIT_OFFSET = 0;
  localparam int REGISTER_3_BIT_FIELD_1_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_3_BIT_FIELD_1_BIT_MASK = 4'hf;
  localparam int REGISTER_3_BIT_FIELD_1_BIT_OFFSET = 4;
  localparam int REGISTER_3_BIT_FIELD_2_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_3_BIT_FIELD_2_BIT_MASK = 4'hf;
  localparam int REGISTER_3_BIT_FIELD_2_BIT_OFFSET = 8;
  localparam int REGISTER_3_BIT_FIELD_3_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_3_BIT_FIELD_3_BIT_MASK = 4'hf;
  localparam int REGISTER_3_BIT_FIELD_3_BIT_OFFSET = 16;
  localparam int REGISTER_4_BYTE_WIDTH = 4;
  localparam int REGISTER_4_BYTE_SIZE = 4;
  localparam bit [7:0] REGISTER_4_BYTE_OFFSET = 8'h0c;
  localparam int REGISTER_4_BIT_FIELD_0_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_4_BIT_FIELD_0_BIT_MASK = 4'hf;
  localparam int REGISTER_4_BIT_FIELD_0_BIT_OFFSET = 0;
  localparam int REGISTER_4_BIT_FIELD_1_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_4_BIT_FIELD_1_BIT_MASK = 4'hf;
  localparam int REGISTER_4_BIT_FIELD_1_BIT_OFFSET = 8;
  localparam int REGISTER_4_BIT_FIELD_2_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_4_BIT_FIELD_2_BIT_MASK = 4'hf;
  localparam int REGISTER_4_BIT_FIELD_2_BIT_OFFSET = 12;
  localparam int REGISTER_4_BIT_FIELD_3_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_4_BIT_FIELD_3_BIT_MASK = 4'hf;
  localparam int REGISTER_4_BIT_FIELD_3_BIT_OFFSET = 16;
  localparam int REGISTER_5_BYTE_WIDTH = 4;
  localparam int REGISTER_5_BYTE_SIZE = 4;
  localparam bit [7:0] REGISTER_5_BYTE_OFFSET = 8'h10;
  localparam int REGISTER_5_BIT_FIELD_0_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_5_BIT_FIELD_0_BIT_MASK = 2'h3;
  localparam int REGISTER_5_BIT_FIELD_0_BIT_OFFSET = 0;
  localparam int REGISTER_5_BIT_FIELD_1_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_5_BIT_FIELD_1_BIT_MASK = 2'h3;
  localparam int REGISTER_5_BIT_FIELD_1_BIT_OFFSET = 2;
  localparam int REGISTER_5_BIT_FIELD_2_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_5_BIT_FIELD_2_BIT_MASK = 2'h3;
  localparam int REGISTER_5_BIT_FIELD_2_BIT_OFFSET = 4;
  localparam int REGISTER_5_BIT_FIELD_3_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_5_BIT_FIELD_3_BIT_MASK = 2'h3;
  localparam int REGISTER_5_BIT_FIELD_3_BIT_OFFSET = 6;
  localparam int REGISTER_5_BIT_FIELD_4_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_5_BIT_FIELD_4_BIT_MASK = 2'h3;
  localparam int REGISTER_5_BIT_FIELD_4_BIT_OFFSET = 8;
  localparam int REGISTER_5_BIT_FIELD_5_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_5_BIT_FIELD_5_BIT_MASK = 2'h3;
  localparam int REGISTER_5_BIT_FIELD_5_BIT_OFFSET = 10;
  localparam int REGISTER_5_BIT_FIELD_6_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_5_BIT_FIELD_6_BIT_MASK = 2'h3;
  localparam int REGISTER_5_BIT_FIELD_6_BIT_OFFSET = 12;
  localparam int REGISTER_5_BIT_FIELD_7_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_5_BIT_FIELD_7_BIT_MASK = 2'h3;
  localparam int REGISTER_5_BIT_FIELD_7_BIT_OFFSET = 14;
  localparam int REGISTER_5_BIT_FIELD_8_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_5_BIT_FIELD_8_BIT_MASK = 2'h3;
  localparam int REGISTER_5_BIT_FIELD_8_BIT_OFFSET = 16;
  localparam int REGISTER_5_BIT_FIELD_9_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_5_BIT_FIELD_9_BIT_MASK = 2'h3;
  localparam int REGISTER_5_BIT_FIELD_9_BIT_OFFSET = 20;
  localparam int REGISTER_5_BIT_FIELD_10_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_5_BIT_FIELD_10_BIT_MASK = 2'h3;
  localparam int REGISTER_5_BIT_FIELD_10_BIT_OFFSET = 22;
  localparam int REGISTER_5_BIT_FIELD_11_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_5_BIT_FIELD_11_BIT_MASK = 2'h3;
  localparam int REGISTER_5_BIT_FIELD_11_BIT_OFFSET = 24;
  localparam int REGISTER_6_BYTE_WIDTH = 8;
  localparam int REGISTER_6_BYTE_SIZE = 8;
  localparam bit [7:0] REGISTER_6_BYTE_OFFSET = 8'h14;
  localparam int REGISTER_6_BIT_FIELD_0_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_6_BIT_FIELD_0_BIT_MASK = 4'hf;
  localparam int REGISTER_6_BIT_FIELD_0_BIT_OFFSET = 0;
  localparam int REGISTER_6_BIT_FIELD_1_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_6_BIT_FIELD_1_BIT_MASK = 4'hf;
  localparam int REGISTER_6_BIT_FIELD_1_BIT_OFFSET = 4;
  localparam int REGISTER_6_BIT_FIELD_2_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_6_BIT_FIELD_2_BIT_MASK = 4'hf;
  localparam int REGISTER_6_BIT_FIELD_2_BIT_OFFSET = 8;
  localparam int REGISTER_6_BIT_FIELD_3_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_6_BIT_FIELD_3_BIT_MASK = 4'hf;
  localparam int REGISTER_6_BIT_FIELD_3_BIT_OFFSET = 12;
  localparam int REGISTER_6_BIT_FIELD_4_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_6_BIT_FIELD_4_BIT_MASK = 4'hf;
  localparam int REGISTER_6_BIT_FIELD_4_BIT_OFFSET = 16;
  localparam int REGISTER_6_BIT_FIELD_5_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_6_BIT_FIELD_5_BIT_MASK = 4'hf;
  localparam int REGISTER_6_BIT_FIELD_5_BIT_OFFSET = 20;
  localparam int REGISTER_6_BIT_FIELD_6_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_6_BIT_FIELD_6_BIT_MASK = 4'hf;
  localparam int REGISTER_6_BIT_FIELD_6_BIT_OFFSET = 24;
  localparam int REGISTER_6_BIT_FIELD_7_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_6_BIT_FIELD_7_BIT_MASK = 4'hf;
  localparam int REGISTER_6_BIT_FIELD_7_BIT_OFFSET = 28;
  localparam int REGISTER_6_BIT_FIELD_8_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_6_BIT_FIELD_8_BIT_MASK = 4'hf;
  localparam int REGISTER_6_BIT_FIELD_8_BIT_OFFSET = 32;
  localparam int REGISTER_6_BIT_FIELD_9_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_6_BIT_FIELD_9_BIT_MASK = 4'hf;
  localparam int REGISTER_6_BIT_FIELD_9_BIT_OFFSET = 36;
  localparam int REGISTER_7_BYTE_WIDTH = 4;
  localparam int REGISTER_7_BYTE_SIZE = 4;
  localparam bit [7:0] REGISTER_7_BYTE_OFFSET = 8'h1c;
  localparam int REGISTER_7_BIT_FIELD_0_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_7_BIT_FIELD_0_BIT_MASK = 4'hf;
  localparam int REGISTER_7_BIT_FIELD_0_BIT_OFFSET = 0;
  localparam int REGISTER_7_BIT_FIELD_1_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_7_BIT_FIELD_1_BIT_MASK = 4'hf;
  localparam int REGISTER_7_BIT_FIELD_1_BIT_OFFSET = 8;
  localparam int REGISTER_7_BIT_FIELD_2_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_7_BIT_FIELD_2_BIT_MASK = 4'hf;
  localparam int REGISTER_7_BIT_FIELD_2_BIT_OFFSET = 16;
  localparam int REGISTER_7_BIT_FIELD_3_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_7_BIT_FIELD_3_BIT_MASK = 4'hf;
  localparam int REGISTER_7_BIT_FIELD_3_BIT_OFFSET = 24;
  localparam int REGISTER_8_BYTE_WIDTH = 8;
  localparam int REGISTER_8_BYTE_SIZE = 8;
  localparam bit [7:0] REGISTER_8_BYTE_OFFSET = 8'h20;
  localparam int REGISTER_8_BIT_FIELD_0_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_8_BIT_FIELD_0_BIT_MASK = 4'hf;
  localparam int REGISTER_8_BIT_FIELD_0_BIT_OFFSET = 0;
  localparam int REGISTER_8_BIT_FIELD_1_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_8_BIT_FIELD_1_BIT_MASK = 4'hf;
  localparam int REGISTER_8_BIT_FIELD_1_BIT_OFFSET = 8;
  localparam int REGISTER_8_BIT_FIELD_2_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_8_BIT_FIELD_2_BIT_MASK = 4'hf;
  localparam int REGISTER_8_BIT_FIELD_2_BIT_OFFSET = 16;
  localparam int REGISTER_8_BIT_FIELD_3_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_8_BIT_FIELD_3_BIT_MASK = 4'hf;
  localparam int REGISTER_8_BIT_FIELD_3_BIT_OFFSET = 24;
  localparam int REGISTER_8_BIT_FIELD_4_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_8_BIT_FIELD_4_BIT_MASK = 4'hf;
  localparam int REGISTER_8_BIT_FIELD_4_BIT_OFFSET = 32;
  localparam int REGISTER_8_BIT_FIELD_5_BIT_WIDTH = 4;
  localparam bit [3:0] REGISTER_8_BIT_FIELD_5_BIT_MASK = 4'hf;
  localparam int REGISTER_8_BIT_FIELD_5_BIT_OFFSET = 40;
  localparam int REGISTER_9_BYTE_WIDTH = 4;
  localparam int REGISTER_9_BYTE_SIZE = 4;
  localparam bit [7:0] REGISTER_9_BYTE_OFFSET = 8'h28;
  localparam int REGISTER_9_BIT_FIELD_0_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_9_BIT_FIELD_0_BIT_MASK = 2'h3;
  localparam int REGISTER_9_BIT_FIELD_0_BIT_OFFSET = 0;
  localparam int REGISTER_9_BIT_FIELD_1_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_9_BIT_FIELD_1_BIT_MASK = 2'h3;
  localparam int REGISTER_9_BIT_FIELD_1_BIT_OFFSET = 2;
  localparam int REGISTER_9_BIT_FIELD_2_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_9_BIT_FIELD_2_BIT_MASK = 2'h3;
  localparam int REGISTER_9_BIT_FIELD_2_BIT_OFFSET = 4;
  localparam int REGISTER_9_BIT_FIELD_3_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_9_BIT_FIELD_3_BIT_MASK = 2'h3;
  localparam int REGISTER_9_BIT_FIELD_3_BIT_OFFSET = 6;
  localparam int REGISTER_9_BIT_FIELD_4_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_9_BIT_FIELD_4_BIT_MASK = 2'h3;
  localparam int REGISTER_9_BIT_FIELD_4_BIT_OFFSET = 8;
  localparam int REGISTER_9_BIT_FIELD_5_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_9_BIT_FIELD_5_BIT_MASK = 2'h3;
  localparam int REGISTER_9_BIT_FIELD_5_BIT_OFFSET = 10;
  localparam int REGISTER_10_BYTE_WIDTH = 4;
  localparam int REGISTER_10_BYTE_SIZE = 32;
  localparam int REGISTER_10_ARRAY_SIZE[1] = '{4};
  localparam bit [7:0] REGISTER_10_BYTE_OFFSET[4] = '{8'h30, 8'h38, 8'h40, 8'h48};
  localparam int REGISTER_10_BIT_FIELD_0_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_10_BIT_FIELD_0_BIT_MASK = 2'h3;
  localparam int REGISTER_10_BIT_FIELD_0_BIT_OFFSET[4] = '{0, 8, 16, 24};
  localparam int REGISTER_10_BIT_FIELD_1_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_10_BIT_FIELD_1_BIT_MASK = 2'h3;
  localparam int REGISTER_10_BIT_FIELD_1_BIT_OFFSET[4] = '{2, 10, 18, 26};
  localparam int REGISTER_10_BIT_FIELD_2_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_10_BIT_FIELD_2_BIT_MASK = 2'h3;
  localparam int REGISTER_10_BIT_FIELD_2_BIT_OFFSET[4] = '{4, 12, 20, 28};
  localparam int REGISTER_11_BYTE_WIDTH = 8;
  localparam int REGISTER_11_BYTE_SIZE = 8;
  localparam int REGISTER_11_ARRAY_SIZE[2] = '{2, 4};
  localparam bit [7:0] REGISTER_11_BYTE_OFFSET[2][4] = '{'{8'h50, 8'h50, 8'h50, 8'h50}, '{8'h50, 8'h50, 8'h50, 8'h50}};
  localparam int REGISTER_11_BIT_FIELD_0_BIT_WIDTH = 8;
  localparam bit [7:0] REGISTER_11_BIT_FIELD_0_BIT_MASK = 8'hff;
  localparam int REGISTER_11_BIT_FIELD_0_BIT_OFFSET[4] = '{0, 16, 32, 48};
  localparam int REGISTER_11_BIT_FIELD_1_BIT_WIDTH = 8;
  localparam bit [7:0] REGISTER_11_BIT_FIELD_1_BIT_MASK = 8'hff;
  localparam int REGISTER_11_BIT_FIELD_1_BIT_OFFSET[4] = '{8, 24, 40, 56};
  localparam int REGISTER_12_BYTE_WIDTH = 8;
  localparam int REGISTER_12_BYTE_SIZE = 8;
  localparam bit [7:0] REGISTER_12_BYTE_OFFSET = 8'h50;
  localparam int REGISTER_12_BIT_FIELD_0_BIT_WIDTH = 1;
  localparam bit REGISTER_12_BIT_FIELD_0_BIT_MASK = 1'h1;
  localparam int REGISTER_12_BIT_FIELD_0_BIT_OFFSET = 0;
  localparam int REGISTER_12_BIT_FIELD_1_BIT_WIDTH = 1;
  localparam bit REGISTER_12_BIT_FIELD_1_BIT_MASK = 1'h1;
  localparam int REGISTER_12_BIT_FIELD_1_BIT_OFFSET = 32;
  localparam int REGISTER_13_BYTE_WIDTH = 4;
  localparam int REGISTER_13_BYTE_SIZE = 4;
  localparam bit [7:0] REGISTER_13_BYTE_OFFSET = 8'h60;
  localparam int REGISTER_13_BIT_FIELD_0_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_13_BIT_FIELD_0_BIT_MASK = 2'h3;
  localparam int REGISTER_13_BIT_FIELD_0_BIT_OFFSET = 0;
  localparam int REGISTER_13_BIT_FIELD_1_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_13_BIT_FIELD_1_BIT_MASK = 2'h3;
  localparam int REGISTER_13_BIT_FIELD_1_BIT_OFFSET = 2;
  localparam int REGISTER_13_BIT_FIELD_2_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_13_BIT_FIELD_2_BIT_MASK = 2'h3;
  localparam int REGISTER_13_BIT_FIELD_2_BIT_OFFSET = 4;
  localparam int REGISTER_13_BIT_FIELD_3_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_13_BIT_FIELD_3_BIT_MASK = 2'h3;
  localparam int REGISTER_13_BIT_FIELD_3_BIT_OFFSET = 6;
  localparam int REGISTER_13_BIT_FIELD_4_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_13_BIT_FIELD_4_BIT_MASK = 2'h3;
  localparam int REGISTER_13_BIT_FIELD_4_BIT_OFFSET = 8;
  localparam int REGISTER_13_BIT_FIELD_5_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_13_BIT_FIELD_5_BIT_MASK = 2'h3;
  localparam int REGISTER_13_BIT_FIELD_5_BIT_OFFSET = 10;
  localparam int REGISTER_13_BIT_FIELD_6_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_13_BIT_FIELD_6_BIT_MASK = 2'h3;
  localparam int REGISTER_13_BIT_FIELD_6_BIT_OFFSET = 12;
  localparam int REGISTER_13_BIT_FIELD_7_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_13_BIT_FIELD_7_BIT_MASK = 2'h3;
  localparam int REGISTER_13_BIT_FIELD_7_BIT_OFFSET = 14;
  localparam int REGISTER_13_BIT_FIELD_8_BIT_WIDTH = 2;
  localparam bit [1:0] REGISTER_13_BIT_FIELD_8_BIT_MASK = 2'h3;
  localparam int REGISTER_13_BIT_FIELD_8_BIT_OFFSET = 16;
  localparam int REGISTER_14_BYTE_WIDTH = 4;
  localparam int REGISTER_14_BYTE_SIZE = 4;
  localparam bit [7:0] REGISTER_14_BYTE_OFFSET = 8'h70;
  localparam int REGISTER_14_BIT_FIELD_0_BIT_WIDTH = 1;
  localparam bit REGISTER_14_BIT_FIELD_0_BIT_MASK = 1'h1;
  localparam int REGISTER_14_BIT_FIELD_0_BIT_OFFSET = 0;
  localparam int REGISTER_15_BYTE_WIDTH = 4;
  localparam int REGISTER_15_BYTE_SIZE = 4;
  localparam bit [7:0] REGISTER_15_BYTE_OFFSET = 8'h74;
  localparam int REGISTER_15_BIT_FIELD_0_BIT_WIDTH = 1;
  localparam bit REGISTER_15_BIT_FIELD_0_BIT_MASK = 1'h1;
  localparam int REGISTER_15_BIT_FIELD_0_BIT_OFFSET = 0;
  localparam int REGISTER_17_BYTE_WIDTH = 4;
  localparam int REGISTER_17_BYTE_SIZE = 128;
  localparam bit [7:0] REGISTER_17_BYTE_OFFSET = 8'h80;
endpackage
