`ifndef UART_CSR_VH
`define UART_CSR_VH
`define UART_CSR_RBR_BIT_WIDTH 8
`define UART_CSR_RBR_BIT_MASK 8'hff
`define UART_CSR_RBR_BIT_OFFSET 0
`define UART_CSR_RBR_BYTE_WIDTH 4
`define UART_CSR_RBR_BYTE_SIZE 4
`define UART_CSR_RBR_BYTE_OFFSET 5'h00
`define UART_CSR_THR_BIT_WIDTH 8
`define UART_CSR_THR_BIT_MASK 8'hff
`define UART_CSR_THR_BIT_OFFSET 0
`define UART_CSR_THR_BYTE_WIDTH 4
`define UART_CSR_THR_BYTE_SIZE 4
`define UART_CSR_THR_BYTE_OFFSET 5'h00
`define UART_CSR_IER_ERBFI_BIT_WIDTH 1
`define UART_CSR_IER_ERBFI_BIT_MASK 1'h1
`define UART_CSR_IER_ERBFI_BIT_OFFSET 0
`define UART_CSR_IER_ETBEI_BIT_WIDTH 1
`define UART_CSR_IER_ETBEI_BIT_MASK 1'h1
`define UART_CSR_IER_ETBEI_BIT_OFFSET 1
`define UART_CSR_IER_ELSI_BIT_WIDTH 1
`define UART_CSR_IER_ELSI_BIT_MASK 1'h1
`define UART_CSR_IER_ELSI_BIT_OFFSET 2
`define UART_CSR_IER_EDSSI_BIT_WIDTH 1
`define UART_CSR_IER_EDSSI_BIT_MASK 1'h1
`define UART_CSR_IER_EDSSI_BIT_OFFSET 3
`define UART_CSR_IER_BYTE_WIDTH 4
`define UART_CSR_IER_BYTE_SIZE 4
`define UART_CSR_IER_BYTE_OFFSET 5'h04
`define UART_CSR_IIR_INTPEND_BIT_WIDTH 1
`define UART_CSR_IIR_INTPEND_BIT_MASK 1'h1
`define UART_CSR_IIR_INTPEND_BIT_OFFSET 0
`define UART_CSR_IIR_INTID2_BIT_WIDTH 3
`define UART_CSR_IIR_INTID2_BIT_MASK 3'h7
`define UART_CSR_IIR_INTID2_BIT_OFFSET 1
`define UART_CSR_IIR_BYTE_WIDTH 4
`define UART_CSR_IIR_BYTE_SIZE 4
`define UART_CSR_IIR_BYTE_OFFSET 5'h08
`define UART_CSR_FCR_FIFOEN_BIT_WIDTH 1
`define UART_CSR_FCR_FIFOEN_BIT_MASK 1'h1
`define UART_CSR_FCR_FIFOEN_BIT_OFFSET 0
`define UART_CSR_FCR_RCVR_FIFO_RESET_BIT_WIDTH 1
`define UART_CSR_FCR_RCVR_FIFO_RESET_BIT_MASK 1'h1
`define UART_CSR_FCR_RCVR_FIFO_RESET_BIT_OFFSET 1
`define UART_CSR_FCR_XMIT_FIFO_RESET_BIT_WIDTH 1
`define UART_CSR_FCR_XMIT_FIFO_RESET_BIT_MASK 1'h1
`define UART_CSR_FCR_XMIT_FIFO_RESET_BIT_OFFSET 2
`define UART_CSR_FCR_DMA_MODE_SELECT_BIT_WIDTH 1
`define UART_CSR_FCR_DMA_MODE_SELECT_BIT_MASK 1'h1
`define UART_CSR_FCR_DMA_MODE_SELECT_BIT_OFFSET 3
`define UART_CSR_FCR_RCVR_FIFO_TRIGGER_LEVEL_BIT_WIDTH 2
`define UART_CSR_FCR_RCVR_FIFO_TRIGGER_LEVEL_BIT_MASK 2'h3
`define UART_CSR_FCR_RCVR_FIFO_TRIGGER_LEVEL_BIT_OFFSET 6
`define UART_CSR_FCR_BYTE_WIDTH 4
`define UART_CSR_FCR_BYTE_SIZE 4
`define UART_CSR_FCR_BYTE_OFFSET 5'h08
`define UART_CSR_LCR_WLS_BIT_WIDTH 2
`define UART_CSR_LCR_WLS_BIT_MASK 2'h3
`define UART_CSR_LCR_WLS_BIT_OFFSET 0
`define UART_CSR_LCR_STB_BIT_WIDTH 1
`define UART_CSR_LCR_STB_BIT_MASK 1'h1
`define UART_CSR_LCR_STB_BIT_OFFSET 2
`define UART_CSR_LCR_PEN_BIT_WIDTH 1
`define UART_CSR_LCR_PEN_BIT_MASK 1'h1
`define UART_CSR_LCR_PEN_BIT_OFFSET 3
`define UART_CSR_LCR_EPS_BIT_WIDTH 1
`define UART_CSR_LCR_EPS_BIT_MASK 1'h1
`define UART_CSR_LCR_EPS_BIT_OFFSET 4
`define UART_CSR_LCR_STICK_PARITY_BIT_WIDTH 1
`define UART_CSR_LCR_STICK_PARITY_BIT_MASK 1'h1
`define UART_CSR_LCR_STICK_PARITY_BIT_OFFSET 5
`define UART_CSR_LCR_SET_BREAK_BIT_WIDTH 1
`define UART_CSR_LCR_SET_BREAK_BIT_MASK 1'h1
`define UART_CSR_LCR_SET_BREAK_BIT_OFFSET 6
`define UART_CSR_LCR_DLAB_BIT_WIDTH 1
`define UART_CSR_LCR_DLAB_BIT_MASK 1'h1
`define UART_CSR_LCR_DLAB_BIT_OFFSET 7
`define UART_CSR_LCR_BYTE_WIDTH 4
`define UART_CSR_LCR_BYTE_SIZE 4
`define UART_CSR_LCR_BYTE_OFFSET 5'h0c
`define UART_CSR_MRC_DTR_BIT_WIDTH 1
`define UART_CSR_MRC_DTR_BIT_MASK 1'h1
`define UART_CSR_MRC_DTR_BIT_OFFSET 0
`define UART_CSR_MRC_RTS_BIT_WIDTH 1
`define UART_CSR_MRC_RTS_BIT_MASK 1'h1
`define UART_CSR_MRC_RTS_BIT_OFFSET 1
`define UART_CSR_MRC_OUT1_BIT_WIDTH 1
`define UART_CSR_MRC_OUT1_BIT_MASK 1'h1
`define UART_CSR_MRC_OUT1_BIT_OFFSET 2
`define UART_CSR_MRC_OUT2_BIT_WIDTH 1
`define UART_CSR_MRC_OUT2_BIT_MASK 1'h1
`define UART_CSR_MRC_OUT2_BIT_OFFSET 3
`define UART_CSR_MRC_LOOP_BACK_BIT_WIDTH 1
`define UART_CSR_MRC_LOOP_BACK_BIT_MASK 1'h1
`define UART_CSR_MRC_LOOP_BACK_BIT_OFFSET 4
`define UART_CSR_MRC_BYTE_WIDTH 4
`define UART_CSR_MRC_BYTE_SIZE 4
`define UART_CSR_MRC_BYTE_OFFSET 5'h10
`define UART_CSR_LSR_DR_BIT_WIDTH 1
`define UART_CSR_LSR_DR_BIT_MASK 1'h1
`define UART_CSR_LSR_DR_BIT_OFFSET 0
`define UART_CSR_LSR_OE_BIT_WIDTH 1
`define UART_CSR_LSR_OE_BIT_MASK 1'h1
`define UART_CSR_LSR_OE_BIT_OFFSET 1
`define UART_CSR_LSR_PE_BIT_WIDTH 1
`define UART_CSR_LSR_PE_BIT_MASK 1'h1
`define UART_CSR_LSR_PE_BIT_OFFSET 2
`define UART_CSR_LSR_FE_BIT_WIDTH 1
`define UART_CSR_LSR_FE_BIT_MASK 1'h1
`define UART_CSR_LSR_FE_BIT_OFFSET 3
`define UART_CSR_LSR_BI_BIT_WIDTH 1
`define UART_CSR_LSR_BI_BIT_MASK 1'h1
`define UART_CSR_LSR_BI_BIT_OFFSET 4
`define UART_CSR_LSR_THRE_BIT_WIDTH 1
`define UART_CSR_LSR_THRE_BIT_MASK 1'h1
`define UART_CSR_LSR_THRE_BIT_OFFSET 5
`define UART_CSR_LSR_TEMT_BIT_WIDTH 1
`define UART_CSR_LSR_TEMT_BIT_MASK 1'h1
`define UART_CSR_LSR_TEMT_BIT_OFFSET 6
`define UART_CSR_LSR_ERROR_IN_RCVR_FIFO_BIT_WIDTH 1
`define UART_CSR_LSR_ERROR_IN_RCVR_FIFO_BIT_MASK 1'h1
`define UART_CSR_LSR_ERROR_IN_RCVR_FIFO_BIT_OFFSET 7
`define UART_CSR_LSR_BYTE_WIDTH 4
`define UART_CSR_LSR_BYTE_SIZE 4
`define UART_CSR_LSR_BYTE_OFFSET 5'h14
`define UART_CSR_MSR_DCTS_BIT_WIDTH 1
`define UART_CSR_MSR_DCTS_BIT_MASK 1'h1
`define UART_CSR_MSR_DCTS_BIT_OFFSET 0
`define UART_CSR_MSR_DDSR_BIT_WIDTH 1
`define UART_CSR_MSR_DDSR_BIT_MASK 1'h1
`define UART_CSR_MSR_DDSR_BIT_OFFSET 1
`define UART_CSR_MSR_TERI_BIT_WIDTH 1
`define UART_CSR_MSR_TERI_BIT_MASK 1'h1
`define UART_CSR_MSR_TERI_BIT_OFFSET 2
`define UART_CSR_MSR_DDCD_BIT_WIDTH 1
`define UART_CSR_MSR_DDCD_BIT_MASK 1'h1
`define UART_CSR_MSR_DDCD_BIT_OFFSET 3
`define UART_CSR_MSR_CTS_BIT_WIDTH 1
`define UART_CSR_MSR_CTS_BIT_MASK 1'h1
`define UART_CSR_MSR_CTS_BIT_OFFSET 4
`define UART_CSR_MSR_DSR_BIT_WIDTH 1
`define UART_CSR_MSR_DSR_BIT_MASK 1'h1
`define UART_CSR_MSR_DSR_BIT_OFFSET 5
`define UART_CSR_MSR_RI_BIT_WIDTH 1
`define UART_CSR_MSR_RI_BIT_MASK 1'h1
`define UART_CSR_MSR_RI_BIT_OFFSET 6
`define UART_CSR_MSR_DCD_BIT_WIDTH 1
`define UART_CSR_MSR_DCD_BIT_MASK 1'h1
`define UART_CSR_MSR_DCD_BIT_OFFSET 7
`define UART_CSR_MSR_BYTE_WIDTH 4
`define UART_CSR_MSR_BYTE_SIZE 4
`define UART_CSR_MSR_BYTE_OFFSET 5'h18
`define UART_CSR_SCRATCH_BIT_WIDTH 8
`define UART_CSR_SCRATCH_BIT_MASK 8'hff
`define UART_CSR_SCRATCH_BIT_OFFSET 0
`define UART_CSR_SCRATCH_BYTE_WIDTH 4
`define UART_CSR_SCRATCH_BYTE_SIZE 4
`define UART_CSR_SCRATCH_BYTE_OFFSET 5'h1c
`define UART_CSR_DLL_BIT_WIDTH 8
`define UART_CSR_DLL_BIT_MASK 8'hff
`define UART_CSR_DLL_BIT_OFFSET 0
`define UART_CSR_DLL_BYTE_WIDTH 4
`define UART_CSR_DLL_BYTE_SIZE 4
`define UART_CSR_DLL_BYTE_OFFSET 5'h00
`define UART_CSR_DLM_BIT_WIDTH 8
`define UART_CSR_DLM_BIT_MASK 8'hff
`define UART_CSR_DLM_BIT_OFFSET 0
`define UART_CSR_DLM_BYTE_WIDTH 4
`define UART_CSR_DLM_BYTE_SIZE 4
`define UART_CSR_DLM_BYTE_OFFSET 5'h04
`endif
